��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��L�+�h�0I��y�������b�~�L�ʬ3�&�;��eW����x�k�Ր�7\�?^ �R����:�{|�h.9��4!�B~����/!���o_mnKD��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m����	-ed%�&ȅ:�SU�� +�"�ж~FPjG�E�\�%m���y$��s%e��i�n�*e���}b��@�'�!�uણ(d��RC�Ѓ���p�4�]8����$�a���#��{��݇(� ��2!_�l?�]��\%Z��0�|���e���d� �a�J��ɯ�z�m�LC�	9��Vo�K(�<��@�(��!g�=����,�W5�z��]�}k�<�q�	�8�*�나s.ײ�U��k���:&��i�^=}��m�aQ�W*z�Z�h���*�HV����P?vb����X.�êPK��fr���U��񆔿�*���~�I���/)Z�$��8��m����(Z(�y:@�@��3��ć~$���p�\��0�=bʖ�C]pMdfg�ۜ{���Du��[w0?e�d�O&4��AѕI]sl;�7��+?�<�_�_P��?C1s�<6�tz9�����o?,����a���T����e�������+��XQ�6bX=���3�K�����	1N6�D��8�YK~�e�`�s��Jt�i��t�MD���y��ʊRU� `�C�h�e6��d�<��a+US��a��t�s�5u�V@�>9nr.P�g�Z��s-���&��"2�� ���6sP���,�J�ٵ�^)��P��S�wXH{��S;��@/.~��J��(����?a�-i�J9縚H��"�W� �S���Қ�=�HʁͰ�?V�����Ɛq�k-�T�d��g	c�4��a!3:YY�� �AQ���k���t����2
��s_�->�`�1��7ɹ�욞�CX��6�3���-X���̤�Y��bя��XQ�P]�� ����V:iK+��֘�\�@������������TTtփ��5���T�94щ�k�f�egY����J
ÄFbgix��i�>䇆&�ƃ�)߃_�H1ښ���32d �:ۘ�����o�ׂ����/������1a*hy�'skѴ���дܧ;��D"R��j'��M<_*˚ErE[�����0�����	���D����S�<n ���X�v(~�u@��m���(b�\��X��u<�6N�dWW��J\$2���x/I%��"U��m`�TG3�*y����/`�����{up���QyF��X8��?���J�:��X�t�a\�[)Y���ԁĀ2�:̢J������r���Ӧ@o���1W�+�#��9��F���û�y7{�'���;�U��#e��qT�N�w(�Ωޖ��v�|i.-������h���M3a=v�sڲ��w�ΐO��1$������&�=�4!���]����2_r���&5-�Tu��ɃC=% Dk��ˁUj�ʪL������ �hr߿n �R#������c��w!�����L0�N�a��w�
�!�Z\;	<�𽐮���(ņ��r�7el����Gl�BE����Vǰ�U,OVҺ�u3�I�Ym3К��0� �z��H�Bz�6�����}��g���2��h��G���_���U�T�^C	�t8˽�oh�2�+�l>���H�`gh'�7���3�ZV��2�耏|N
T�f~{��?�����lԜH2 �:�&��V{{������^��jM%�~�	�)@���4��]�i���nr��w�3�Y��@@M{tOLC������í%�
7��uO�	2������Cp�b��P�e��(�v�r*y�I�
JVRh&-[_�Q�z*�,�n7myo&�c�� C�d�'ߍۘ$�'C��2�bӞ�c Ë�h������>Wݪ�4��捯�eD�Q��c�H�qs�"���
�㵙�Xt�d�bH̡uv*�"�>�d�d�x&q�h3�/������/�0@'�"b��x_�0:�Jb�T����������o�80�\Xl�����!
��A$;��	���6�O#C�
	d������q��YwiD;V~�q�w�yl�_�Ė�b��{ʈ%��U�\�t�5��M�~mNk��������3�s�?��׫���*SZ%'j�=����`JLH�aE�6˩g�G@ĉ��-,��h��l猪F������l!�xk�0���UK��I1�n�)NoLPM���h�.�=�(�A_upsʦL�Q8�bxn�?�>竣��R�X-<d���e�Ůe�F�q��Y˷�������i�{?��$�a�գKV�lN��[A�����N��b��w~˝ ҆q��^63���,��2C��D��M�R�?��#v9j �a%��� �Hk��wl�oDY3ӽ�r�ܦ������|C�}�BNC�T`�߲�3��� ��~i�k��Bʠ��]�^V5��yY��,j��>˄�FA��~��:�z
"�[n7.�JR�!����ѡDD����_�0ii疎gz�j���9󽓵��c�i�G(8�K|���ʯ犚��+�?��:��-C"JD9Z��.�o�j,����3P͕	(@;A�=�_��]�M_������]���oq�Q$a�̓C��A�1r�[��&Sd=D�����0&��G
ĩ\�v�]�]�2���Np�!�$����KX�qNY�<���)������8��r�
B>�lJ����W�I���MT~�1�*�~ƛ���Uu ��i}?�fWmñ�Eu}Z�D �}��]��Jz��w�����T��u!8��1	 ��ҩĀb��`{�܉����CC�
�L*��>q�n�T����?4�h�X�?^���^D+z�fc�P\u��N� k��?���I�
�@�:3%J�a�L���J�ʽ#1�(V�ж����7��E���w���<Xc[�=$�\�V��e�{�C!����#�*�t�,#2Wd�=�������#�z R�'��vk��0���i��Y�HX@Oख�-���4��a�9��怅(j��P�E����q��/( <�n��
N����t�TXCmx�e�%YG!�)������kg���'n$������y���k�_�bʉ�Kwi��p�_(P�ab�l�[
���\J�����QP|�E�M7����W����R� s�=����q׬�O�T�N���i��K��>_�h��5)T�|���hUP�t�H; ��)��`�7{4�B�M�mq|Q�j�0'�sm`/�(�n�m`͟p^�^�� �d��Z��a�����W�?\\��I��x|b�'��C�F�%۲�'lK����B33��Hú�Ԧ|`]�P�y2,-����^�6*�xim;d��>�I���/N+S~?D�-L �Q���pu���u���`�>�:�B�ޟ�l��*$N}Q�+���_xZ����<��61[juQL`�9����@��K��e`�$JLਃ�+P�����YT�9��1���ς���?X�@�d���Ɔ|J�ѼÍ�a$r��,�t�yY�=��㺍�JE>{�b[|e2��Is�h��x�G*?ĳz_?��)W�,��t��;�����1C��D��Λr؈�CTE��H�T��:N7����I@-Fa�k�(�̨���0F
�Eq� أ}��b:-ܔ���p~l�@YC��y3 �;|=y|�>���P��a��ū!h72u���>p�0�W5�E4D#_�\4��ֺ�C���H�g>��k!|�DG/]D�lkFh�?�?N�1�6���_�%�o���|���#}��x��.�� &|k/7f�9�d���8ߟ�u�D�c@�Z�]+�������'��!�g������9���M�d��̶�����$�@z�ߝ�9�{��(G\��N�֗f�H�@%X���F�[f�3����9w�B�=a�2��?	�������;h�����.��M�=1k�|1���E�Pp�6�b ��s�1�H6�a@4���I�8-��p:g	���fdK=�,�7ir󷓉�4��-?��Y�r�^xg����y�!-pv^���U�Ёn����b#'���/���Dws�$���m��g��{l+������F�C���N�Sx���̚�P�@����d�uAhr���k��(��'�]��[M��?�����u;���,D��eB��lN	[\/ڑ�٢v��_]j�S����KE��0�F䒫�2����f�lW1z�v�`�P��6�p��}>�%cZQ�	�μ�j�����p�8��oQe}H-Hk��o>����xvQ�(YA0.��]~|-�B|#��0���{� =p3�I���%�����L�;���Z~�=��՞���YF��&�Q^xO�1}l27y��q��d�F�cT���g�:3�)s�U�PA�E��C��l������3/��.�ϝ+�42�@ba"�7�eo���7fAp6��( �!�k�� -�5�: �?bY��WB�X8��q+%7��<^���O�b�4��w����6V'n�dX�_�<K��d���	�:��-�:W�y3%���45���E��7�)��21������oZ&j�?\��</H���\���}��>@q7�fv̹7��"8��=
l���|�9�ݖhg�2iގ�O(����?���=t.�ւ[ľ�f*����@���6]Ѩt��(���	��°U��AW
F��8g�MQ]�V�������Ā�j�ї����$oS�GΞ���{��o"����b!N�P��un&����Z>.��<�a�=%��#]צ�6?���G+[�WJ/v�~(a�:�V���g�B&H����#��ھ�߳�Fҷ|�A�NX�?�G��t=]� Ǯ�����r\#�rg�E��O<��k�Pr���Z[���������7$�>T���,is�����ԴB��0�����1�^�#J���`�ƹ9cgV8���L�1`. �;v%W"�D� W��y将ݩ�+6��]~�sa�*Q҅���a+<�LZ���ɗ�_l������Gl~{������X@������K(#���ӏ>�d����Mʜc��]>_�/�
'�n�ik����o� ���)���vw��`�Bh�Lb.F'�p}�D�D"ǉ��o[X�Ү[�7�{�`^�t��r�����y���^"��Re�!X���M�p �g��4�������¶�𾠇�fD�u��g�9��QvF�:��;�7�ˀ��v�;�\���ή����8�خ!f��fNڞ�d
`;g������S��>��[�����_yA[�ɢ�E��7���k=p7M���	y_c�h�2���ƚ?��#ɭ��h��$���7}�G���5K�M�Q�{)B}�u�UN��b�F� �ֺxh��'H9�k�e9�t�ZX���jI�|�S߷�k�hW��VZ����ʵ���ȳu��� ���ɥ�G4���S��6ɪ�!�¾l(�P�G}��*���~gny*F��)�#�Ҭ�I���)t�H-,�HSb.��R��Z濸ja:���	.�>����e���K"�Hk��/�\>�śQ�i�:�!�]�q#������W�ʢ�_\�ao��?�O!���?����"*k�.]���֎���r�����ufB���2WvK��{!N�)���h��]Κ�!A��p�(mL-{� �����MB�o���zZ�t��Ϧ����1k#��MP3a7�`2_�O�uǭc�)\G��-���X7�k���&MmrZ���fێދ�%�~��EPI�E{�`�|0z�b�I#=j��j���(g�8���m��C�q������#".��3�ٻ�����B�֓�6����S1�>C#X����a�?u+C��V����2gBm���H��:�5H�8q�����0��T�p�ub��p�1L<�3�(���zC&��#AB��W�@���N(�)7��G헻h�+�D��f5����\M�ϖ�9΁h�+p]��^�i��!x7����K�C��2�~��-�O�&@Ş��/�~QrU�~��/%50Y1�"2p"�F|q���3XL_���իT��0^� aw�o��4u�ƣ���rqI=Z6\VG`3jǲ����m���?�7���w��a�/��px��a�N�q�;n/�56��S���\��<�df#J�9�[��M\Q�.F�҄0�.谻����7�	7�9�F�1ŧ��!��!��}rRUhrf�p�2E�~QQ�j�dgw�q�ـ\}`�g{fc+jo�m��W"�� ���b$o`A��"�}���7�H֔��:cV��SA���ά�������9�ݍ�g@���R>ڳVO9dh�e�s�rgj�W�Ҩ巂*6жg{Q��xP�	FMz�����U^���Jn�����#H�j4B08����$�)��QsBp⊛l�@�|���tnS����@l�j��)�r�Y_+��Y�i97��(7�I�y(+r�g����z�%%��^";�:�G���ѡ�V}�Q�b�Ǣi;Į4�$�~����B�vz����a��,�2�jA':��ˬ]]Ș\�Ś�{��=�q��,.���1��rH�s������˚adQ�5��N��J\�#Nbk��9�\��}.f~��O̶=3��cA4������
=Q��[e�dy�Ch���M9A�E3�t[����8�P�8��Um�n���@�r��b�&�]��� L=�~Lu�5kJ��n�Z�+� �V�%k�i��{�6x�V�D����_Eg� `�|
��vf��mE��mrR�w��nP���Z��ҫ�RF}��;��f{��/y��+|Ȩ�h�� ����p�h\������:JI�s0z���Q4�:L4ԗ�+�δ�G�~�c���V��6b��B�F�[�@*�)������t��2dV�ޟ��|ʌ�֮��Y����h��Y^?8�����M�<���Jq�����;��6z�_?6W�Z�E��H�Ѓ{����ET`WF�7�b!#�6vy��D�>F��F	�L	�}���Y*h\:��)Wds�i����X�%�k�^����V��Z�E�}m��g
ra�}"���s=�Ip��IK{9��h�z{q>�Ĵ�Sݶ|�Mi��J(��#���8���T'��!����u俚ݜR)�炨s���m��T|
��V4At<��4;\OV%1d`^.�<�����Yދ'���7l���۲Z40�g��ym5P�pͯ4�pA�_-�4E$�V �-���'F���Z�LF��!kB�P~��{�������M	�q�������u��מKj`�3ce����ڞ1���,����(�2�OS:�ӜlV_C	��\ZptULU��Ƈr�-}r<�&�&\����s�)̢��B;4|6A�B�c�$P��Q��T����-(޼$��W�mex
�9u̲�f�x�P���̽�gC�Z��	2O�<�:�a�DL\����O���#hs�����M�!�{lz������[c���aM�ڀ�ۏ���26|q��I����6��y�Y�m�|�A�rX&^2},6��Z �t1�J)I*�e�(ƀ�҄&��֘�x�H�>��?M��ؕ�2g��c��B��(��h.���4�0�yn�z�IǢq��mNA�����X��ҳ��se6���γ��戥^14��	��H���y��1�i����pR<���\m��@����V	�)1����Pߐ����C|��4E.�Nm�Wr�5��E��b���	�4!����Z�<��Hs��y=>N�u�I �W�ی�)u/���:S����We		�%&K��`MA)Nx�S�Y\�S�M�	��x�b�1�"��#B=u�����mE��%��p
�<���b܇u��|8��-�����s���%��`����m�/�=�C�89[�+)�Z���A�W��٫����c,���
��)�-�Vw��epJZƥ����q������t�ׂ��L�d��5kp�2QJȘ�w����?��3�?��R��*L���`�g�q:Յ�K�n��;ގȍE����� �-������B�f#�G(TC��M����Hu>0��_��)��^x�3z6�x�M�����Q���{�@���r���]%�����r�R�����[���������`@v�"� ;�[�e��i���2��W��s�zk�G�\*�pi�� Z�N�@?x�`<���5B�.N��^��@Ԯ֯��N�H'h���{o٨N��PT��>�����3����ꢵ�,�����g�� s�U��/�����Ay��B�N�?l��W�ZKp�� h�t����\��!��w:�{(�tu�`;�A@R�Iő6��]y�N��(q��e���! �5k�㐠$���w*D�����=�w��gS3���x,�Է#�Q71%c���*o�@qk�
�&��WA?������ӑu��x�cm.G���ˇNܠr+h���"T[��ߝ�׽�=�Gqf����p^"�t�9�#��n�C�8�/��p	#}�@ր&�_��'��	#��@op����C�A^ޮ��w&�}�H����T�N+���� ��2�i��X�7����k�γ)y?4uD�^���mk�F����@�(֋�gY�W�S���^�c��^F� ��gE�7D�E]�W�̨O��cc��%�����ǚ��R�0���e�F����wG�lV6�wL�S�ƸT�?m�W�r�����u�������ӄ[��2y��oj�T
8��y	�u	;��N��)u�ОT��M�T�X4Xyn����ʨq��ֻ������b�N�%`�i����xi��JW]՛��ƒ���U�,�3*���D�9�wfa,�;Z�1���ؤ���8Q=��/�lz<�����ϥn�|�Me�&���p��Ne���|�ޚ�LT�J�7�wy8�y:N(1<ܾN��2N�ka<����I+q�aQ�ת(#yh�Z��U_e��K���K��C@Ix�2��}u|��)�݊��c��|v�l�X���qe�9��gJ�J���~����(�(���dk2Il��b��R.u2�9Xe1#�q���/Ύ�@�ϫ�f�B��6�T�>�`ɚ�5�IL͓��q�*�ygj���E4C[����d��\�u3=�UIql7�/�9�y#I�o_�^q�=I�Ώ²lj�������ܑ�V�/�	�1J]�� ��0'��ϲ�@z| ڏ ����S����LW��_�#z;�h[,`��~��c��c|y/F5��ǉ�d��bu#�r�E�T�jd��������·HG�5 C~��6�"`�|&t�ӈ�D��{��
ZDW�}��$d��G�v$��Ư��|�/��>��� kʶ��-��0��TP��kZ_m���GK�'&Q�$v�~w�0#��p��brSj�,3.���eI��aR��H���R��]���o$��S�8=�SA�ȈK������ 5��5��\:0��+��E:4�i��h�?��z#���u�@�RG`*=E�))�+D�+��Y�#�22�*��*��m&CTA��?���}�֔������(�h���	ܦ���a���XXK�敃��DH��|��n��H-����z�[)*���	!@׫�|����V�����!�b��}6j;��������J8�Ս�r��t��d���"Q����*�qf*�� X���Th?2y�S���v��6�<���˃ý�Q.z��U��E^�ڇ'Q�aG���`��������6�t�B�Z)��F�	�Hޚ
��s�%�Y|�ӊ�Ou�kpG"��,4I L��K?�M���H�JX��"1��0�k\����_^ ��r�'�K�n�������5�H�S�;�Q�j�H�.w���u����U�=P�ۖ�<`x�	OJ� ��:���zLk.D=W���ӕb�ݣ������V͊IxP}-�����nTl���-a'��4�ab����u������D��,������y�Z[dUu�]�¯�I��ܕ�	N����V��w�v��J��o������߈Oo���n��M�涍=��5䞛*ș]� 솎�7c\/�����@d�G=���z��V�+���,�L�=��o��G$:�I/ě7L#�_-�~�~*mD��E�s����]Ϧ5�ydλ�'ن�����D+�	�ޯ�E�n ��e���8@�^��ܺ�n��L�B ܐ��K�U-��,����ѣ�����$u~�o�����1���������^��(pG�ك��.̗���e���C� tV���2���k�*p�F�tY	����~��ج�V�� t4�ƒ�Qd�-��G���x���w�Vռ����z�.�N�0�D�[|X���D��*B��]��5�C�K�ODô��b��ܠ�	%��h�	�L�[���w�;���~f�d�U���ǛG?�Sک���d���� ��ͯ�8m�oբ�?n����<7�����u>1��,:��EJ
7OoP$f9@���럭_�Id U
v�#�?Ff��=�L���Y����%�!�붚�hR�l5� ����*iw�sa������`p�;n�$�P\�JIXڼ�u(UK��󭕺Bs$,�i3�+k���4���N�	�⹿��:��0�`�/�������J�����Q�dG��d)R�G*E#㓌������`��%&�$ԛt��������>+.��V�y��Nl> {i0��I�sU��PQ�C��}+�@�zݡ�[Jԩ��g�Z�T�]|D��v���d� J>?�xt<ܑ܌iG��+L���	,��s։���~��4�+��)��;"n_�q�ŗ�|rA�͆�����ST�h��OD���΋��ECe& ��P�:zH`"Kf[(�3_��x�p�����Ŗ\��`Ɗ[I�Sc�9u9��Lw8�J�:�),�=���Ve�2ޥt�5�ъ�1$OKp(���pح-�y����z�Uf�Ȋp�8.WC�e�W,+v��m����9��p]lzo0$0��g�I�>��Vi�����m�WÐ���`��g^�^5jE�/���:��?e�_)���{?v�Z��b��.U~h*ry�NH�?���)�)��\c�6�D�_���|ₛ�ω��a5�G��P�D9�n��_9k=�B��(i������Tb�Ml�߉$	8f�-n�72���IBՐu��\Ew��9Bt?��8�YGKhP��:~����`N��Pss�N��9�ȭ��M�z��Pb�Tc�s����G�P��O��X@�K�(�ϙ